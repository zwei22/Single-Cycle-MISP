module SIGN_EXT(
    in,
    out
);

input   [15:0] in;
output  [31:0] out;

assign out = in;

endmodule